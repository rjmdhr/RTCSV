`timescale 1ns/1ns

module rtc_driver_tb;

    logic clk;
    logic [2:0] push_but;
    logic rst;
    logic man_sw;
    logic [5:0] sev_seg[6:0];

    // tb driver/check logic
    logic [] test_vec [1000:0]
    logic 

    rtc_driver UUT (
        .
    )


endmodule