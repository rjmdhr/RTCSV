`timescale 1ns/100ps

// This module takes a reference clock and drives 6 7-segment displays to display
// the time in HH:MM:SS format. It also contains a toggle switch for a time set mode
// and 3 push buttons to set the time columns. The accuracy will be limited to the
// internal clock
// DE2-115 SOC board
// note: switches are default logic 0 when in "down position"
//       buttons are active low (logic high when not pressed)
module rtc_driver(
	input logic clk, //50 MHz clock (20ns)
	input logic [2:0] push_but, //increase digit
	input logic rst, // master reset
	input logic man_sw, //manual clock set
	output logic [5:0] sev_seg[7:0] //6 displays, arranged in pin format;
	// 10-9-1-2-4-6-7 | g-f-e-d-c-b-a.

	// total input|outputs = 6|48
);

// divisors for 1Hz and 1kHz clock enables
parameter div1kHz = 24999; //50E6/25E3 = 2000x ~/sec
parameter div1Hz = 24999999; //50E6/25E6 = 2x ~/sec

logic [24:0] cnt1Hz;
logic cnten; //count enable
logic [15:0] cnt1kHz;
logic shiften; //shift reg enable

// counters (1 is 10s column, 0 is 1s column)
logic [3:0] sec1, sec0;
logic [3:0] min1, min0;
logic [1:0] hr1, hr0;

//seven segment output registers
//0 for 1s column, 1 for 10s column
logic [6:0] ssH0, ssH1, ssM0, ssM1, ssS0, ssS1;

/** 1Hz clock enable for displays */
always_ff @(posedge clk or negedge rst) begin
	if (rst == 1'b0) begin
		cnt1Hz <= 25'd0;
		cnten <= 1'b0;
	end
	else begin
		if (cnt1Hz == div1Hz) begin
			cnten <= 1'b1;
			cnt1Hz <= 25'd0;
		end
		else begin
			cnten <= 1'b0;
			cnt1Hz <= cnt1Hz + 25'd1;
		end
	end
end

/** 1kHz clock enable for shift register debouncers */
always_ff @(posedge clk or negedge rst) begin
	if (rst == 1'b0) begin
		cnt1kHz <= 16'd0;
		shiftten <= 1'b0;
	end
	else begin
		if (cnt1Hz == div1kHz) begin
			shiften <= 1'b1;
			cnt1kHz <= 16'd0;
		end
		else begin
			shiften <= 1'b0;
			cnt1kHz <= cnt1kHz + 16'd1;
		end
	end
end

/* Button debouncers */
always_ff @(posedge clk50M or negedge resetn) begin
	
end

/** HH:MM:SS counters */
// seconds counter - increments and resets at 59
always_ff @(posedge clk50M or negedge resetn) begin : seconds_counter
	if (resetn == 1'b0) begin
		sec0 <= 4'd0;
		sec1 <= 4'd0;
	end
	else begin
		// auto
		if (~man_switch) begin
			if (count_en) begin
				if (sec0 < 4'd9) begin
					sec0 <= sec0 + 4'd1;
				end
				else begin
					if (sec1 == 4'd5) begin
						sec1 <= 4'd0;
						sec0 <= 4'd0;
					end
					else begin
						sec1 <= sec1 + 4'd1;
						sec0 <= 4'd0;
					end
				end
			end
		end
		// manual
		else begin
			
		end
	end
end
// minutes counter - increments every minute at the seconds reset
always_ff @(posedge clk50M or negedge resetn) begin : minutes_counter
	if (resetn == 1'b0) begin
		min_ctr_0 <= 4'd0;
		min_ctr_1 <= 4'd0;
	end
	else begin
		// auto
		if (~man_switch) begin
			if (count_en) begin
				if (sec1 == 4'd5 && sec0 == 4'd9) begin
					if (min_ctr_0 < 4'd9) begin
						min_ctr_0 <= min_ctr_0 + 4'd1;
					end
					else begin
						if (min_ctr_1 == 4'd5) begin
							min_ctr_1 <= 4'd0;
							min_ctr_0 <= 4'd0;
						end
						else begin
							min_ctr_1 <= min_ctr_1 + 4'd1;
							min_ctr_0 <= 4'd0;
						end
					end
				end
			end
		end
		// manual
		else begin
			
		end
	end
end
// hours counter - increments every hour at the seconds reset (24 hour time)
always_ff @(posedge clk50M or negedge resetn) begin : hours_counter
	if (resetn == 1'b0) begin
		hr_ctr_0 <= 4'd0;
		hr_ctr_1 <= 4'd0;
	end
	else begin
		// auto
		if (~man_switch) begin
			if (count_en) begin
				if (sec1 == 4'd5 && sec0 == 4'd9) begin
					if (min_ctr_1 == 4'd5 && min_ctr_0 == 4'd9) begin
						if (hr_ctr_1 == 2'd2 && hr_ctr_0 == 4'd3) begin
							hr_ctr_1 <= 2'd0;
							hr_ctr_0 <= 4'd0;
						end
						else begin
							if (hr_ctr_0 < 4'd9) begin
								hr_ctr_0 <= hr_ctr_0 + 4'd1;
							end
							else begin
								hr_ctr_1 <= hr_ctr_1 + 2'd1;
								hr_ctr_0 <= 4'd0;
							end
						end
					end
				end
			end
		end
		// manual
		else begin
			
		end
	end
end

endmodule